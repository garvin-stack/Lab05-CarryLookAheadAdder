//=========================================================================
// Name & Email must be EXACTLY as in Gradescope roster!
// Name: 
// Email: 
// 
// Assignment name: 
// Lab section: 
// TA: 
// 
// I hereby certify that I have not received assistance on this assignment,
// or used code, from ANY outside source other than the instruction team
// (apart from what was provided in the starter file).
//
//=========================================================================

`timescale 1ns / 1ps

//  Constant definitions 

module carry_look_ahead_logic # (parameter NUMBITS = 4) (
    input  wire [NUMBITS-1:0] p, 
    input  wire [NUMBITS-1:0] g,
    input  wire c_in,
    output reg  [NUMBITS:0] c
);

    // ------------------------------
    // Insert your solution below
    // ------------------------------ 

endmodule